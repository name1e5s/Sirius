`timescale 1ns / 1ps
// Dual issue detect engine.
module dual_engine(
        input                           alpha_issue,
        input [31:0]                    instruction_alpha,
        input [31:0]                    instruction_beta,
        output logic                    beta_issue
);

// TODO：

endmodule